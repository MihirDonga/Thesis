
// testbench_pkg.sv
`ifndef TESTBENCH_PKG_SV
`define TESTBENCH_PKG_SV
package testbench_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "uart_cov_pkg.sv"
  `include "apb_cov_pkg.sv"

  // UART
  `include "uart_config.sv"
  `include "apb_config.sv"
  `include "uart_transaction.sv"
  `include "apb_transaction.sv"
  `include "uart_sequencer.sv"
  `include "apb_sequencer.sv"
  `include "uart_sequence.sv"
  `include "apb_sequence.sv"
  `include "uart_driver.sv"
  `include "apb_driver.sv"
  `include "uart_monitor.sv"
  `include "apb_monitor.sv"
  `include "uart_agent.sv"
  `include "apb_agent.sv"

  // Virtual Sequencer & Sequences
  `include "apbuart_vsequencer.sv"
  `include "apbuart_vseq_base.sv"


  // Scoreboard
  `include "apbuart_scoreboard.sv"

  // Tests
  `include "apbuart_environment.sv"
  `include "apbuart_base_test.sv"
  `include "apbuart_config_test.sv"
  `include "apbuart_data_compare_test.sv"
  `include "apbuart_frame_error_test.sv"
  `include "apbuart_free_error_test.sv"
  `include "apbuart_parity_error_test.sv"
  `include "apbuart_rec_drv_test.sv"
  `include "apbuart_rec_readreg_test.sv"


endpackage : testbench_pkg

`endif